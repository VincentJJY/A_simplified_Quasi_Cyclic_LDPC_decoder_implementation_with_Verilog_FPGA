`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2024/05/19 23:46:54
// Design Name: 
// Module Name: VariableNodeProcessingUnit_tb
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module VariableNodeProcessingUnit_tb;

    // Testbench signals
    reg clk;
    reg rst;
    reg [15:0] I1;
    reg [15:0] I2;
    reg [15:0] I3;
    reg [15:0] I4;
    reg [15:0] Z;
    wire [15:0] L1;
    wire [15:0] L2;
    wire [15:0] L3;
    wire [15:0] L4;
    wire C;

    // Instantiate the DUT (Device Under Test)
    VariableNodeProcessingUnit dut (
        .clk(clk),
        .rst(rst),
        .I1(I1),
        .I2(I2),
        .I3(I3),
        .I4(I4),
        .Z(Z),
        .L1(L1),
        .L2(L2),
        .L3(L3),
        .L4(L4),
        .C(C)
    );

    initial clk=0;
    always #10 clk = ~clk;


    initial begin
        rst = 1;
        I1  = 16'b0;
        I2  = 16'b0;
        I3  = 16'b0;
        I4  = 16'b0;
        Z   = 16'b0;
        #10;
        @(posedge clk) rst = 0;
        #10;
        I1 = 16'b000101;         
        I2 = 16'b001010; 
        I3 = 16'b001111; 
        I4 = 16'b010100; 
        Z  = 16'b000011; 
        #20;
        I1 = 16'b111011; 
        I2 = 16'b111010; 
        I3 = 16'b111001; 
        I4 = 16'b111000; 
        Z  = 16'b111110;  
        #20;
        I1 = 16'b010101; 
        I2 = 16'b011010; 
        I3 = 16'b011111; 
        I4 = 16'b100100; 
        Z  = 16'b000111;  

        #20;
        I1 = 16'b1101100111011010; 
        I2 = 16'b0111101111101010; 
        I3 = 16'b0001101000110001; 
        I4 = 16'b1101100010101011; 
        Z = 16'b1110001010100010; 
        #20;

        I1 = 16'b0111101101001110; 
        I2 = 16'b1000010101011100; 
        I3 = 16'b0101110001011100; 
        I4 = 16'b0101000011101101; 
        Z = 16'b0000000011000100; 
        #20;

        I1 = 16'b1000001110001000; 
        I2 = 16'b1110101010011011; 
        I3 = 16'b0000111110110111; 
        I4 = 16'b1100001000000100; 
        Z = 16'b1100001011000001; 
        #20;

        I1 = 16'b0010110100111001; 
        I2 = 16'b1001011100010101; 
        I3 = 16'b0111101001101111; 
        I4 = 16'b1100100011100100; 
        Z = 16'b1011101111100100; 
        #20;

        I1 = 16'b0011001011000100; 
        I2 = 16'b0000110100110101; 
        I3 = 16'b1111001001110001; 
        I4 = 16'b0110000010010010; 
        Z = 16'b1110101110100000; 
        #20;

        I1 = 16'b0010111000110111; 
        I2 = 16'b1001100000010111; 
        I3 = 16'b1101011000110110; 
        I4 = 16'b1010000101000100; 
        Z = 16'b0101010100011101; 
        #20;

        I1 = 16'b1111010010011010; 
        I2 = 16'b1101111000110111; 
        I3 = 16'b1111000000011111; 
        I4 = 16'b0010111001110010; 
        Z = 16'b0100101011000000; 
        #20;

        I1 = 16'b1010101100110101; 
        I2 = 16'b1011111000111010; 
        I3 = 16'b0010000011111111; 
        I4 = 16'b0111101001111101; 
        Z = 16'b0111111111001010; 
        #20;

        I1 = 16'b1101000000000101; 
        I2 = 16'b1010001100110010; 
        I3 = 16'b0001101110111111; 
        I4 = 16'b0000100001011100; 
        Z = 16'b0010101111000110; 
        #20;

        I1 = 16'b0001000110101110; 
        I2 = 16'b1000100000100000; 
        I3 = 16'b1000001110011101; 
        I4 = 16'b0010011111101100; 
        Z = 16'b1011001011100011; 
        #20;

        I1 = 16'b1010010111101110; 
        I2 = 16'b0011100010010100; 
        I3 = 16'b1000100001011011; 
        I4 = 16'b0101001010001001; 
        Z = 16'b0011000001110100; 
        #20;

        I1 = 16'b0000000011100011; 
        I2 = 16'b1001100001010100; 
        I3 = 16'b0110101110000011; 
        I4 = 16'b0000001110011110; 
        Z = 16'b1000100111101110; 
        #20;

        I1 = 16'b1101010000011101; 
        I2 = 16'b1100100111100101; 
        I3 = 16'b1111100110101100; 
        I4 = 16'b0001011101010001; 
        Z = 16'b0010101011110111; 
        #20;

        I1 = 16'b0000110101101011; 
        I2 = 16'b1111000001100111; 
        I3 = 16'b1101001101111110; 
        I4 = 16'b1101010000011101; 
        Z = 16'b1100110010100111; 
        #20;

        I1 = 16'b0000010011000011; 
        I2 = 16'b1000101101001111; 
        I3 = 16'b0101110110111010; 
        I4 = 16'b1001101110010011; 
        Z = 16'b1100001101010101; 
        #20;

        I1 = 16'b1010010101110110; 
        I2 = 16'b0110000000001010; 
        I3 = 16'b0011111000011110; 
        I4 = 16'b1101111001011100; 
        Z = 16'b0011100101101111; 
        #20;

        I1 = 16'b1111001101110111; 
        I2 = 16'b1010011101011100; 
        I3 = 16'b0111110100111011; 
        I4 = 16'b0001011001111001; 
        Z = 16'b1101000100001100; 
        #20;

        I1 = 16'b1111010000000100; 
        I2 = 16'b1111111000010010; 
        I3 = 16'b1111001111110001; 
        I4 = 16'b1110110110110001; 
        Z = 16'b1011110010001010; 
        #20;

        I1 = 16'b1101011000001111; 
        I2 = 16'b0101010111110011; 
        I3 = 16'b1011011011011110; 
        I4 = 16'b0110000010000000; 
        Z = 16'b0000010100000000; 
        #20;

        I1 = 16'b0011100010000010; 
        I2 = 16'b1101111010011001; 
        I3 = 16'b1110101011000001; 
        I4 = 16'b0100001111000001; 
        Z = 16'b1100111111010000; 
        #20;

        I1 = 16'b1010010110011100; 
        I2 = 16'b1111101001011000; 
        I3 = 16'b1000000001011001; 
        I4 = 16'b0010111101011100; 
        Z = 16'b0111101101001011; 
        #20;

        I1 = 16'b1111001000111001; 
        I2 = 16'b1100111010100011; 
        I3 = 16'b0001100011001001; 
        I4 = 16'b0111011010001101; 
        Z = 16'b0110101001100101; 
        #20;

        I1 = 16'b1100111110100011; 
        I2 = 16'b1111100011110110; 
        I3 = 16'b1000010000010001; 
        I4 = 16'b0110110110011101; 
        Z = 16'b1110000001100000; 
        #20;

        I1 = 16'b0101000001011100; 
        I2 = 16'b0110011011010011; 
        I3 = 16'b0111000100110001; 
        I4 = 16'b0010110011110100; 
        Z = 16'b0111101011100111; 
        #20;

        I1 = 16'b1111010010010000; 
        I2 = 16'b0100001011110010; 
        I3 = 16'b1110100011110101; 
        I4 = 16'b1111001000011101; 
        Z = 16'b1110101110100110; 
        #20;

        I1 = 16'b1100000101010110; 
        I2 = 16'b0000011101011011; 
        I3 = 16'b1110001100111011; 
        I4 = 16'b0001101100111100; 
        Z = 16'b1110111011011010; 
        #20;

        I1 = 16'b1001000011001011; 
        I2 = 16'b1101111101100101; 
        I3 = 16'b1110011111101101; 
        I4 = 16'b1010000010001011; 
        Z = 16'b1011000101110010; 
        #20;

        I1 = 16'b0001111000110001; 
        I2 = 16'b1000101011111010; 
        I3 = 16'b0010111101110111; 
        I4 = 16'b0001110111001110; 
        Z = 16'b0110001111011000; 
        #20;

        I1 = 16'b0111101000010111; 
        I2 = 16'b0111010010001001; 
        I3 = 16'b0111010101011000; 
        I4 = 16'b1101100010000111; 
        Z = 16'b1101000110010110; 
        #20;

        I1 = 16'b0111010110010010; 
        I2 = 16'b1111101011100111; 
        I3 = 16'b1000000100000100; 
        I4 = 16'b0011010111010011; 
        Z = 16'b0110100010010111; 
        #20;

        I1 = 16'b1001101111110010; 
        I2 = 16'b1010010110010000; 
        I3 = 16'b0100010100011011; 
        I4 = 16'b1110000100010011; 
        Z = 16'b0001010110101100; 
        #20;

        I1 = 16'b1100101101110011; 
        I2 = 16'b1101111010111111; 
        I3 = 16'b0000000110010011; 
        I4 = 16'b0110010001100101; 
        Z = 16'b0000001011110011; 
        
        #90;

        
        $stop;
    end

    // Monitor signals
    initial begin
        $monitor("Time=%0d, rst=%b, I1=%b, I2=%b, I3=%b, I4=%b, Z=%b, L1=%b, L2=%b, L3=%b, L4=%b, C=%b",
                 $time, rst, I1, I2, I3, I4, Z, L1, L2, L3, L4, C);
    end
endmodule
