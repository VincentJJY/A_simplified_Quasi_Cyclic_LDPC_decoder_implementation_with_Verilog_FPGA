`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2024/05/19 18:24:59
// Design Name: 
// Module Name: CheckNodeProcessingUnit_tb
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////
// delay : 5 cycles

module CheckNodeProcessingUnit_tb;

// Inputs
reg clk;
reg rst;
reg [15:0] Lcn_0;
reg [15:0] Lcn_1;
reg [15:0] Lcn_2;
reg [15:0] Lcn_3;
reg [15:0] Lcn_4;
reg [15:0] Lcn_5;
reg [15:0] Lcn_6;
reg [15:0] Lcn_7;
reg [15:0] Lcn_8;
reg [15:0] Lcn_9;
reg [15:0] Lcn_10;
reg [15:0] Lcn_11;
reg [15:0] Lcn_12;
reg [15:0] Lcn_13;
reg [15:0] Lcn_14;
reg [15:0] Lcn_15;
reg [15:0] Lcn_16;
reg [15:0] Lcn_17;
reg [15:0] Lcn_18;
reg [15:0] Lcn_19;
reg [15:0] Lcn_20;
reg [15:0] Lcn_21;
reg [15:0] Lcn_22;
reg [15:0] Lcn_23;
reg [15:0] Lcn_24;
reg [15:0] Lcn_25;
reg [15:0] Lcn_26;
reg [15:0] Lcn_27;
reg [15:0] Lcn_28;
reg [15:0] Lcn_29;
reg [15:0] Lcn_30;
reg [15:0] Lcn_31;
wire [15:0] sign_magnitude_0 ; 
wire [15:0] sign_magnitude_1 ; 
wire [15:0] sign_magnitude_2 ; 
wire [15:0] sign_magnitude_3 ;
wire [15:0] sign_magnitude_4 ; 
wire [15:0] sign_magnitude_5 ; 
wire [15:0] sign_magnitude_6 ; 
wire [15:0] sign_magnitude_7 ;
wire [15:0] sign_magnitude_8 ; 
wire [15:0] sign_magnitude_9 ; 
wire [15:0] sign_magnitude_10; 
wire [15:0] sign_magnitude_11;
wire [15:0] sign_magnitude_12; 
wire [15:0] sign_magnitude_13; 
wire [15:0] sign_magnitude_14; 
wire [15:0] sign_magnitude_15;
wire [15:0] sign_magnitude_16; 
wire [15:0] sign_magnitude_17; 
wire [15:0] sign_magnitude_18; 
wire [15:0] sign_magnitude_19;
wire [15:0] sign_magnitude_20; 
wire [15:0] sign_magnitude_21; 
wire [15:0] sign_magnitude_22; 
wire [15:0] sign_magnitude_23;
wire [15:0] sign_magnitude_24; 
wire [15:0] sign_magnitude_25; 
wire [15:0] sign_magnitude_26; 
wire [15:0] sign_magnitude_27;
wire [15:0] sign_magnitude_28; 
wire [15:0] sign_magnitude_29; 
wire [15:0] sign_magnitude_30; 
wire [15:0] sign_magnitude_31; 



// Instantiate the Unit Under Test (UUT)
CheckNodeProcessingUnit uut (
    .clk(clk), 
    .rst(rst), 
    .Lcn_0(Lcn_0), 
    .Lcn_1(Lcn_1), 
    .Lcn_2(Lcn_2), 
    .Lcn_3(Lcn_3), 
    .Lcn_4(Lcn_4), 
    .Lcn_5(Lcn_5), 
    .Lcn_6(Lcn_6), 
    .Lcn_7(Lcn_7), 
    .Lcn_8(Lcn_8), 
    .Lcn_9(Lcn_9), 
    .Lcn_10(Lcn_10), 
    .Lcn_11(Lcn_11), 
    .Lcn_12(Lcn_12), 
    .Lcn_13(Lcn_13), 
    .Lcn_14(Lcn_14), 
    .Lcn_15(Lcn_15), 
    .Lcn_16(Lcn_16), 
    .Lcn_17(Lcn_17), 
    .Lcn_18(Lcn_18), 
    .Lcn_19(Lcn_19), 
    .Lcn_20(Lcn_20), 
    .Lcn_21(Lcn_21), 
    .Lcn_22(Lcn_22), 
    .Lcn_23(Lcn_23), 
    .Lcn_24(Lcn_24), 
    .Lcn_25(Lcn_25), 
    .Lcn_26(Lcn_26), 
    .Lcn_27(Lcn_27), 
    .Lcn_28(Lcn_28), 
    .Lcn_29(Lcn_29), 
    .Lcn_30(Lcn_30), 
    .Lcn_31(Lcn_31), 
    .sign_magnitude_0 (  sign_magnitude_0  ), 
    .sign_magnitude_1 (  sign_magnitude_1  ), 
    .sign_magnitude_2 (  sign_magnitude_2  ), 
    .sign_magnitude_3 (  sign_magnitude_3  ),
    .sign_magnitude_4 (  sign_magnitude_4  ), 
    .sign_magnitude_5 (  sign_magnitude_5  ), 
    .sign_magnitude_6 (  sign_magnitude_6  ), 
    .sign_magnitude_7 (  sign_magnitude_7  ),
    .sign_magnitude_8 (  sign_magnitude_8  ), 
    .sign_magnitude_9 (  sign_magnitude_9  ), 
    .sign_magnitude_10(  sign_magnitude_10 ), 
    .sign_magnitude_11(  sign_magnitude_11 ),
    .sign_magnitude_12(  sign_magnitude_12 ), 
    .sign_magnitude_13(  sign_magnitude_13 ), 
    .sign_magnitude_14(  sign_magnitude_14 ), 
    .sign_magnitude_15(  sign_magnitude_15 ),
    .sign_magnitude_16(  sign_magnitude_16 ), 
    .sign_magnitude_17(  sign_magnitude_17 ), 
    .sign_magnitude_18(  sign_magnitude_18 ), 
    .sign_magnitude_19(  sign_magnitude_19 ),
    .sign_magnitude_20(  sign_magnitude_20 ), 
    .sign_magnitude_21(  sign_magnitude_21 ), 
    .sign_magnitude_22(  sign_magnitude_22 ), 
    .sign_magnitude_23(  sign_magnitude_23 ),
    .sign_magnitude_24(  sign_magnitude_24 ), 
    .sign_magnitude_25(  sign_magnitude_25 ), 
    .sign_magnitude_26(  sign_magnitude_26 ), 
    .sign_magnitude_27(  sign_magnitude_27 ),
    .sign_magnitude_28(  sign_magnitude_28 ), 
    .sign_magnitude_29(  sign_magnitude_29 ), 
    .sign_magnitude_30(  sign_magnitude_30 ), 
    .sign_magnitude_31(  sign_magnitude_31 )  
);

initial  clk=0     ;
always #10 clk = ~clk;


initial begin

    rst = 1;
    Lcn_0 = 0;
    Lcn_1 = 0;
    Lcn_2 = 0;
    Lcn_3 = 0;
    Lcn_4 = 0;
    Lcn_5 = 0;
    Lcn_6 = 0;
    Lcn_7 = 0;
    Lcn_8 = 0;
    Lcn_9 = 0;
    Lcn_10 = 0;
    Lcn_11 = 0;
    Lcn_12 = 0;
    Lcn_13 = 0;
    Lcn_14 = 0;
    Lcn_15 = 0;
    Lcn_16 = 0;
    Lcn_17 = 0;
    Lcn_18 = 0;
    Lcn_19 = 0;
    Lcn_20 = 0;
    Lcn_21 = 0;
    Lcn_22 = 0;
    Lcn_23 = 0;
    Lcn_24 = 0;
    Lcn_25 = 0;
    Lcn_26 = 0;
    Lcn_27 = 0;
    Lcn_28 = 0;
    Lcn_29 = 0;
    Lcn_30 = 0;
    Lcn_31 = 0;


    #20;
    @(posedge clk) rst = 0;
    #20;
    

    Lcn_0  = 16'b000001;
    Lcn_1  = 16'b000010;
    Lcn_2  = 16'b000011;
    Lcn_3  = 16'b000100;
    Lcn_4  = 16'b000101;
    Lcn_5  = 16'b000110;
    Lcn_6  = 16'b000111;
    Lcn_7  = 16'b001000;
    Lcn_8  = 16'b001001;
    Lcn_9  = 16'b001010;
    Lcn_10 = 16'b001011;
    Lcn_11 = 16'b001100;
    Lcn_12 = 16'b001101;
    Lcn_13 = 16'b001110;
    Lcn_14 = 16'b001111;
    Lcn_15 = 16'b010000;
    Lcn_16 = 16'b010001;
    Lcn_17 = 16'b010010;
    Lcn_18 = 16'b010011;
    Lcn_19 = 16'b010100;
    Lcn_20 = 16'b010101;
    Lcn_21 = 16'b010110;
    Lcn_22 = 16'b010111;
    Lcn_23 = 16'b011000;
    Lcn_24 = 16'b011001;
    Lcn_25 = 16'b011010;
    Lcn_26 = 16'b011011;
    Lcn_27 = 16'b011100;
    Lcn_28 = 16'b011101;
    Lcn_29 = 16'b011110;
    Lcn_30 = 16'b011111;
    Lcn_31 = 16'b100000;
    #20;


    Lcn_0  = 16'b111111;
    Lcn_1  = 16'b111110;
    Lcn_2  = 16'b111101;
    Lcn_3  = 16'b111100;
    Lcn_4  = 16'b111011;
    Lcn_5  = 16'b111010;
    Lcn_6  = 16'b111001;
    Lcn_7  = 16'b111000;
    Lcn_8  = 16'b110111;
    Lcn_9  = 16'b110110;
    Lcn_10 = 16'b110101;
    Lcn_11 = 16'b110100;
    Lcn_12 = 16'b110011;
    Lcn_13 = 16'b110010;
    Lcn_14 = 16'b110001;
    Lcn_15 = 16'b110000;
    Lcn_16 = 16'b101111;
    Lcn_17 = 16'b101110;
    Lcn_18 = 16'b101101;
    Lcn_19 = 16'b101100;
    Lcn_20 = 16'b101011;
    Lcn_21 = 16'b101010;
    Lcn_22 = 16'b101001;
    Lcn_23 = 16'b101000;
    Lcn_24 = 16'b100111;
    Lcn_25 = 16'b100110;
    Lcn_26 = 16'b100101;
    Lcn_27 = 16'b100100;
    Lcn_28 = 16'b100011;
    Lcn_29 = 16'b100010;
    Lcn_30 = 16'b100001;
    Lcn_31 = 16'b100000;
    #20;


    Lcn_0  = 16'b101001;
    Lcn_1  = 16'b010110;
    Lcn_2  = 16'b001001;
    Lcn_3  = 16'b111000;
    Lcn_4  = 16'b000100;
    Lcn_5  = 16'b011101;
    Lcn_6  = 16'b101110;
    Lcn_7  = 16'b010001;
    Lcn_8  = 16'b110000;
    Lcn_9  = 16'b001100;
    Lcn_10 = 16'b111101;
    Lcn_11 = 16'b100010;
    Lcn_12 = 16'b011011;
    Lcn_13 = 16'b000111;
    Lcn_14 = 16'b101100;
    Lcn_15 = 16'b010011;
    Lcn_16 = 16'b110100;
    Lcn_17 = 16'b001111;
    Lcn_18 = 16'b111010;
    Lcn_19 = 16'b100101;
    Lcn_20 = 16'b011000;
    Lcn_21 = 16'b000001;
    Lcn_22 = 16'b101011;
    Lcn_23 = 16'b010101;
    Lcn_24 = 16'b110001;
    Lcn_25 = 16'b001011;
    Lcn_26 = 16'b111110;
    Lcn_27 = 16'b100100;
    Lcn_28 = 16'b011010;
    Lcn_29 = 16'b000010;
    Lcn_30 = 16'b101111;
    Lcn_31 = 16'b010100;

    #20;
    Lcn_0 = 16'b0011000011111000;
    Lcn_1 = 16'b1011100111111100;
    Lcn_2 = 16'b0101011110101101;
    Lcn_3 = 16'b0010110011001001;
    Lcn_4 = 16'b1000111100001000;
    Lcn_5 = 16'b1110101010101110;
    Lcn_6 = 16'b0111110011111111;
    Lcn_7 = 16'b1111101110111001;
    Lcn_8 = 16'b1100001010011010;
    Lcn_9 = 16'b0010010001000010;
    Lcn_10 = 16'b1010010010101100;
    Lcn_11 = 16'b0101111000011000;
    Lcn_12 = 16'b0000011000000000;
    Lcn_13 = 16'b0111100101111101;
    Lcn_14 = 16'b0101000001011010;
    Lcn_15 = 16'b0001100100100100;
    Lcn_16 = 16'b1101000100110111;
    Lcn_17 = 16'b0100110000010010;
    Lcn_18 = 16'b0010110010000011;
    Lcn_19 = 16'b1000001010001111;
    Lcn_20 = 16'b0111010101010011;
    Lcn_21 = 16'b0000000100010011;
    Lcn_22 = 16'b1011001100010001;
    Lcn_23 = 16'b1011010111001100;
    Lcn_24 = 16'b0100100100111011;
    Lcn_25 = 16'b0000011101010110;
    Lcn_26 = 16'b0000100111001110;
    Lcn_27 = 16'b0110111101101100;
    Lcn_28 = 16'b1001100110100100;
    Lcn_29 = 16'b1111101000101011;
    Lcn_30 = 16'b1100111100101101;
    Lcn_31 = 16'b1000000101010110;
    
    #20;
    Lcn_0 = 16'b1111000100000011;
    Lcn_1 = 16'b1111100101101001;
    Lcn_2 = 16'b0010100111010000;
    Lcn_3 = 16'b1001100110010010;
    Lcn_4 = 16'b0001001001110101;
    Lcn_5 = 16'b1111110010110100;
    Lcn_6 = 16'b1100000101110111;
    Lcn_7 = 16'b0011011111111110;
    Lcn_8 = 16'b1110011010001110;
    Lcn_9 = 16'b0111110000001010;
    Lcn_10 = 16'b1001000101001100;
    Lcn_11 = 16'b1111001100001110;
    Lcn_12 = 16'b0101001011001111;
    Lcn_13 = 16'b1101010001110101;
    Lcn_14 = 16'b0111110011110011;
    Lcn_15 = 16'b0111101010000100;
    Lcn_16 = 16'b0001011010111000;
    Lcn_17 = 16'b0000101001100100;
    Lcn_18 = 16'b1001001100110010;
    Lcn_19 = 16'b1000101000100110;
    Lcn_20 = 16'b0001101010101111;
    Lcn_21 = 16'b1000011011110011;
    Lcn_22 = 16'b1101111000001000;
    Lcn_23 = 16'b0100110001010010;
    Lcn_24 = 16'b1001110001101110;
    Lcn_25 = 16'b1000100110110000;
    Lcn_26 = 16'b1001101111011000;
    Lcn_27 = 16'b0110000010101100;
    Lcn_28 = 16'b0100010100110000;
    Lcn_29 = 16'b0100101111101011;
    Lcn_30 = 16'b1010001111000100;
    Lcn_31 = 16'b0010111101100011;
    
    #20;
    Lcn_0 = 16'b0101000101111000;
    Lcn_1 = 16'b0011000010010011;
    Lcn_2 = 16'b0100011110100010;
    Lcn_3 = 16'b1110000000011110;
    Lcn_4 = 16'b1010111000001110;
    Lcn_5 = 16'b0011100000111110;
    Lcn_6 = 16'b0111111100000000;
    Lcn_7 = 16'b0101001010001110;
    Lcn_8 = 16'b1000100001111100;
    Lcn_9 = 16'b1000001001000011;
    Lcn_10 = 16'b1011101001111001;
    Lcn_11 = 16'b0011101011100011;
    Lcn_12 = 16'b1001011100100110;
    Lcn_13 = 16'b0100000100001110;
    Lcn_14 = 16'b0010011010001100;
    Lcn_15 = 16'b1111100011100001;
    Lcn_16 = 16'b0100110011111110;
    Lcn_17 = 16'b1101011100111010;
    Lcn_18 = 16'b1101100001010001;
    Lcn_19 = 16'b1111110001011010;
    Lcn_20 = 16'b1001101101010011;
    Lcn_21 = 16'b0100111111111111;
    Lcn_22 = 16'b0111110110011011;
    Lcn_23 = 16'b1010110001010011;
    Lcn_24 = 16'b0101101111011000;
    Lcn_25 = 16'b1101101110010000;
    Lcn_26 = 16'b1011010011010011;
    Lcn_27 = 16'b1110010000100111;
    Lcn_28 = 16'b1101100001011111;
    Lcn_29 = 16'b1000110001010101;
    Lcn_30 = 16'b0010010100010001;
    Lcn_31 = 16'b0011101011111110;
    
    #20;
    Lcn_0 = 16'b0100011111011010;
    Lcn_1 = 16'b0000101110011111;
    Lcn_2 = 16'b0110110011000101;
    Lcn_3 = 16'b0001001011011011;
    Lcn_4 = 16'b1000110010011111;
    Lcn_5 = 16'b1101101101101000;
    Lcn_6 = 16'b1010011101001101;
    Lcn_7 = 16'b1001010111100110;
    Lcn_8 = 16'b1101010010001110;
    Lcn_9 = 16'b1010101111000011;
    Lcn_10 = 16'b1110101000100110;
    Lcn_11 = 16'b0101001111010001;
    Lcn_12 = 16'b1110111110111111;
    Lcn_13 = 16'b0100100111001010;
    Lcn_14 = 16'b1101111110010010;
    Lcn_15 = 16'b1000110010101011;
    Lcn_16 = 16'b1001110101100011;
    Lcn_17 = 16'b0111110110000101;
    Lcn_18 = 16'b1110111101101010;
    Lcn_19 = 16'b1111111100000011;
    Lcn_20 = 16'b0001000111001000;
    Lcn_21 = 16'b0101011100001110;
    Lcn_22 = 16'b1110110100110001;
    Lcn_23 = 16'b0101110000001000;
    Lcn_24 = 16'b0010111000111001;
    Lcn_25 = 16'b1101000001000010;
    Lcn_26 = 16'b0110111010101100;
    Lcn_27 = 16'b1011110111011010;
    Lcn_28 = 16'b1100000000111010;
    Lcn_29 = 16'b0011100100101100;
    Lcn_30 = 16'b0001110011101111;
    Lcn_31 = 16'b1001100111011011;
    
    #20;
    Lcn_0 = 16'b0111100001011010;
    Lcn_1 = 16'b1000010110011101;
    Lcn_2 = 16'b1010000001000011;
    Lcn_3 = 16'b0001101001010111;
    Lcn_4 = 16'b1001010011111001;
    Lcn_5 = 16'b0111100101000110;
    Lcn_6 = 16'b0000011101100100;
    Lcn_7 = 16'b0001100110010010;
    Lcn_8 = 16'b0000110100100000;
    Lcn_9 = 16'b0001100101100001;
    Lcn_10 = 16'b1001111100110100;
    Lcn_11 = 16'b0010100000010110;
    Lcn_12 = 16'b0100110000111010;
    Lcn_13 = 16'b1011111111010011;
    Lcn_14 = 16'b0100111011100111;
    Lcn_15 = 16'b1001101001000100;
    Lcn_16 = 16'b1111001001101001;
    Lcn_17 = 16'b1001100100111101;
    Lcn_18 = 16'b1101000101100101;
    Lcn_19 = 16'b0010000001111010;
    Lcn_20 = 16'b1011100111010011;
    Lcn_21 = 16'b0110100100011001;
    Lcn_22 = 16'b0001000110011001;
    Lcn_23 = 16'b1000001111000010;
    Lcn_24 = 16'b0100001101000110;
    Lcn_25 = 16'b0010000001010100;
    Lcn_26 = 16'b0100100101110010;
    Lcn_27 = 16'b0011001100011010;
    Lcn_28 = 16'b0011011000000101;
    Lcn_29 = 16'b0100000100110111;
    Lcn_30 = 16'b1110101000110011;
    Lcn_31 = 16'b0000011110011110;
    
    #20;
    Lcn_0 = 16'b0011100000001100;
    Lcn_1 = 16'b0011010110010001;
    Lcn_2 = 16'b1001001100010110;
    Lcn_3 = 16'b0111110010011011;
    Lcn_4 = 16'b0010101111110110;
    Lcn_5 = 16'b1100100101100100;
    Lcn_6 = 16'b0110011011100100;
    Lcn_7 = 16'b1111011100101101;
    Lcn_8 = 16'b1101001101000001;
    Lcn_9 = 16'b0001101100010000;
    Lcn_10 = 16'b0110110010001111;
    Lcn_11 = 16'b1010100000000110;
    Lcn_12 = 16'b0101001101000110;
    Lcn_13 = 16'b0011010010110000;
    Lcn_14 = 16'b0101100110111010;
    Lcn_15 = 16'b0101010000100011;
    Lcn_16 = 16'b0001010101000010;
    Lcn_17 = 16'b1101001101011100;
    Lcn_18 = 16'b1111010101100110;
    Lcn_19 = 16'b1110011101110110;
    Lcn_20 = 16'b1101110011010100;
    Lcn_21 = 16'b1010110100100100;
    Lcn_22 = 16'b0101011100110100;
    Lcn_23 = 16'b0100010101110010;
    Lcn_24 = 16'b0011111000111110;
    Lcn_25 = 16'b1111000010101001;
    Lcn_26 = 16'b0011100000001011;
    Lcn_27 = 16'b1000110110101011;
    Lcn_28 = 16'b0000001010000011;
    Lcn_29 = 16'b0111000011000010;
    Lcn_30 = 16'b1101001101100010;
    Lcn_31 = 16'b1111111011101001;
    
    #20;
    Lcn_0 = 16'b0010010101101001;
    Lcn_1 = 16'b1010110011110111;
    Lcn_2 = 16'b0101110100110000;
    Lcn_3 = 16'b1101111100011011;
    Lcn_4 = 16'b1111000010110111;
    Lcn_5 = 16'b0001110110010100;
    Lcn_6 = 16'b1110100101010001;
    Lcn_7 = 16'b1111110101100000;
    Lcn_8 = 16'b1010010011100111;
    Lcn_9 = 16'b1111111000001011;
    Lcn_10 = 16'b0101011001001100;
    Lcn_11 = 16'b0011001110101100;
    Lcn_12 = 16'b1110000111100100;
    Lcn_13 = 16'b0010010000011110;
    Lcn_14 = 16'b0001001000010101;
    Lcn_15 = 16'b0100110011000100;
    Lcn_16 = 16'b1001010110100111;
    Lcn_17 = 16'b0100110101111011;
    Lcn_18 = 16'b0001011110111010;
    Lcn_19 = 16'b0111101011010100;
    Lcn_20 = 16'b0001000101110011;
    Lcn_21 = 16'b1001011100001101;
    Lcn_22 = 16'b0100110001010000;
    Lcn_23 = 16'b0110111110100010;
    Lcn_24 = 16'b1100100111101000;
    Lcn_25 = 16'b0111100011101011;
    Lcn_26 = 16'b0111101110111000;
    Lcn_27 = 16'b1111000001001011;
    Lcn_28 = 16'b0111011110000111;
    Lcn_29 = 16'b1110001101000000;
    Lcn_30 = 16'b1001111010000110;
    Lcn_31 = 16'b1000110100001100;
    
    #20;
    Lcn_0 = 16'b1010111110111010;
    Lcn_1 = 16'b0100110111111010;
    Lcn_2 = 16'b0010010101010001;
    Lcn_3 = 16'b0010001000001100;
    Lcn_4 = 16'b0101000011000110;
    Lcn_5 = 16'b1011010001110010;
    Lcn_6 = 16'b0011010111101101;
    Lcn_7 = 16'b0011001000010001;
    Lcn_8 = 16'b1101101100001010;
    Lcn_9 = 16'b1111010010010100;
    Lcn_10 = 16'b0010111001010000;
    Lcn_11 = 16'b1100010011011100;
    Lcn_12 = 16'b1101101011110110;
    Lcn_13 = 16'b1011011110011101;
    Lcn_14 = 16'b1111011101110111;
    Lcn_15 = 16'b0000010111100001;
    Lcn_16 = 16'b0100010001101011;
    Lcn_17 = 16'b0111011110001110;
    Lcn_18 = 16'b1010110101011011;
    Lcn_19 = 16'b1000011100001010;
    Lcn_20 = 16'b1010000111100100;
    Lcn_21 = 16'b1000110010110001;
    Lcn_22 = 16'b0100101100110010;
    Lcn_23 = 16'b0000011111001011;
    Lcn_24 = 16'b1101111010100011;
    Lcn_25 = 16'b1101010110000100;
    Lcn_26 = 16'b0110110111101101;
    Lcn_27 = 16'b1111110110010111;
    Lcn_28 = 16'b1101101001110011;
    Lcn_29 = 16'b1011100001011010;
    Lcn_30 = 16'b0001111111100001;
    Lcn_31 = 16'b1001100011000110;
    
    #20;
    Lcn_0 = 16'b0101110111100010;
    Lcn_1 = 16'b1100011001100111;
    Lcn_2 = 16'b0100111100001000;
    Lcn_3 = 16'b0101101000001101;
    Lcn_4 = 16'b1100110111101110;
    Lcn_5 = 16'b1101000101100101;
    Lcn_6 = 16'b0100010101010100;
    Lcn_7 = 16'b0010111001110110;
    Lcn_8 = 16'b1110110010101000;
    Lcn_9 = 16'b1110100101110011;
    Lcn_10 = 16'b1110111110110110;
    Lcn_11 = 16'b1000101100101001;
    Lcn_12 = 16'b1011110010101110;
    Lcn_13 = 16'b0110111100010101;
    Lcn_14 = 16'b0000010010111110;
    Lcn_15 = 16'b1101101010101100;
    Lcn_16 = 16'b1001100111111111;
    Lcn_17 = 16'b0111000111011101;
    Lcn_18 = 16'b1001100101111100;
    Lcn_19 = 16'b1111001111111010;
    Lcn_20 = 16'b1101110001100111;
    Lcn_21 = 16'b0011110111110001;
    Lcn_22 = 16'b1101111010010000;
    Lcn_23 = 16'b0101100010100101;
    Lcn_24 = 16'b0100010100111010;
    Lcn_25 = 16'b0011100100111100;
    Lcn_26 = 16'b0011101101100100;
    Lcn_27 = 16'b0010011111011011;
    Lcn_28 = 16'b0101011111001100;
    Lcn_29 = 16'b0101110100100111;
    Lcn_30 = 16'b0101111011111000;
    Lcn_31 = 16'b0000010011110010;
    
    #20;
    Lcn_0 = 16'b0001111011010101;
    Lcn_1 = 16'b1011010111010110;
    Lcn_2 = 16'b1000101001001000;
    Lcn_3 = 16'b0010010100001011;
    Lcn_4 = 16'b1100010110001010;
    Lcn_5 = 16'b0001111100001110;
    Lcn_6 = 16'b1111111111000110;
    Lcn_7 = 16'b1110001000111001;
    Lcn_8 = 16'b0101101000000001;
    Lcn_9 = 16'b0001100101111111;
    Lcn_10 = 16'b1111010101111101;
    Lcn_11 = 16'b1100001110100010;
    Lcn_12 = 16'b0101100011001010;
    Lcn_13 = 16'b0101111110010100;
    Lcn_14 = 16'b0001101100100011;
    Lcn_15 = 16'b1011110000010000;
    Lcn_16 = 16'b1001011000010011;
    Lcn_17 = 16'b1110110011011010;
    Lcn_18 = 16'b0110001110000010;
    Lcn_19 = 16'b0000110010011111;
    Lcn_20 = 16'b0001111001101011;
    Lcn_21 = 16'b1110100101010110;
    Lcn_22 = 16'b1001110010101001;
    Lcn_23 = 16'b0011000010111110;
    Lcn_24 = 16'b0011100011110010;
    Lcn_25 = 16'b0011011111011010;
    Lcn_26 = 16'b0111010101010101;
    Lcn_27 = 16'b0011111110001010;
    Lcn_28 = 16'b1101011011100111;
    Lcn_29 = 16'b1100111000111110;
    Lcn_30 = 16'b0011101000000001;
    Lcn_31 = 16'b0100010001010100;
    
    #20;
    Lcn_0 = 16'b0101101000100100;
    Lcn_1 = 16'b1000000110100100;
    Lcn_2 = 16'b0010011001010110;
    Lcn_3 = 16'b0110011010001011;
    Lcn_4 = 16'b1010010010010010;
    Lcn_5 = 16'b1000101100011000;
    Lcn_6 = 16'b0111000100001010;
    Lcn_7 = 16'b1100010100010000;
    Lcn_8 = 16'b0101011110001000;
    Lcn_9 = 16'b0001000111100001;
    Lcn_10 = 16'b1111000000011000;
    Lcn_11 = 16'b0110100011010110;
    Lcn_12 = 16'b0000011011100000;
    Lcn_13 = 16'b0100011100001001;
    Lcn_14 = 16'b0101000111100110;
    Lcn_15 = 16'b1111000100010110;
    Lcn_16 = 16'b1010011110100000;
    Lcn_17 = 16'b0011001100010110;
    Lcn_18 = 16'b0001101110001000;
    Lcn_19 = 16'b1101011001110111;
    Lcn_20 = 16'b0001110011011111;
    Lcn_21 = 16'b0101011100011010;
    Lcn_22 = 16'b0100010111110011;
    Lcn_23 = 16'b0100000110000011;
    Lcn_24 = 16'b0011000110011000;
    Lcn_25 = 16'b1110101010111110;
    Lcn_26 = 16'b1011011010100111;
    Lcn_27 = 16'b1100100010110101;
    Lcn_28 = 16'b0010010111111010;
    Lcn_29 = 16'b1000100100011011;
    Lcn_30 = 16'b0010110010010110;
    Lcn_31 = 16'b1011101010001011;
    
    #20;
    Lcn_0 = 16'b1011011100011101;
    Lcn_1 = 16'b1010000100111010;
    Lcn_2 = 16'b0010110111111100;
    Lcn_3 = 16'b0010010011000000;
    Lcn_4 = 16'b1001110011011001;
    Lcn_5 = 16'b1011111000010110;
    Lcn_6 = 16'b0110001111011011;
    Lcn_7 = 16'b0100110101010011;
    Lcn_8 = 16'b1110101001010110;
    Lcn_9 = 16'b0111011000111111;
    Lcn_10 = 16'b0000110001000010;
    Lcn_11 = 16'b1111001011100001;
    Lcn_12 = 16'b0111001011010011;
    Lcn_13 = 16'b0000111010110011;
    Lcn_14 = 16'b1011110101010010;
    Lcn_15 = 16'b0011010011100001;
    Lcn_16 = 16'b1000011010011011;
    Lcn_17 = 16'b0101111000100101;
    Lcn_18 = 16'b1010001100101111;
    Lcn_19 = 16'b0111101001100001;
    Lcn_20 = 16'b1000011000100101;
    Lcn_21 = 16'b1010101011011001;
    Lcn_22 = 16'b0001100011011100;
    Lcn_23 = 16'b0110101101101010;
    Lcn_24 = 16'b0010010100110100;
    Lcn_25 = 16'b1011101110111100;
    Lcn_26 = 16'b0100000110101010;
    Lcn_27 = 16'b1101111111101100;
    Lcn_28 = 16'b1100101000100100;
    Lcn_29 = 16'b0010010111011111;
    Lcn_30 = 16'b1010100000001011;
    Lcn_31 = 16'b0101010011000000;
    
    #20;
    Lcn_0 = 16'b1110000010110011;
    Lcn_1 = 16'b1000011100111011;
    Lcn_2 = 16'b0111101001110010;
    Lcn_3 = 16'b0111001100001010;
    Lcn_4 = 16'b1010000011010011;
    Lcn_5 = 16'b1100110001001010;
    Lcn_6 = 16'b1011000101011100;
    Lcn_7 = 16'b1011111001101010;
    Lcn_8 = 16'b0111001000010010;
    Lcn_9 = 16'b1110111010100000;
    Lcn_10 = 16'b1001110011101000;
    Lcn_11 = 16'b0111100001000101;
    Lcn_12 = 16'b0110101110100100;
    Lcn_13 = 16'b1111100110100110;
    Lcn_14 = 16'b1010111101110010;
    Lcn_15 = 16'b0010010001100000;
    Lcn_16 = 16'b1000011000100001;
    Lcn_17 = 16'b0010101010100000;
    Lcn_18 = 16'b0011111001001001;
    Lcn_19 = 16'b0111010101001001;
    Lcn_20 = 16'b1011110010111110;
    Lcn_21 = 16'b0000111001111111;
    Lcn_22 = 16'b0000000001000000;
    Lcn_23 = 16'b0101001101110001;
    Lcn_24 = 16'b0110011100000011;
    Lcn_25 = 16'b0101101111000111;
    Lcn_26 = 16'b1001001110000010;
    Lcn_27 = 16'b1000110010110001;
    Lcn_28 = 16'b0101001011100010;
    Lcn_29 = 16'b0101001100100010;
    Lcn_30 = 16'b1101000111000001;
    Lcn_31 = 16'b1000001011010100;
    
    #20;
    Lcn_0 = 16'b0110110000101010;
    Lcn_1 = 16'b0000111100000011;
    Lcn_2 = 16'b0010100001100000;
    Lcn_3 = 16'b1011101101100110;
    Lcn_4 = 16'b0010011110001001;
    Lcn_5 = 16'b0011101101000010;
    Lcn_6 = 16'b1011000011010010;
    Lcn_7 = 16'b0001011001011010;
    Lcn_8 = 16'b1110100101100011;
    Lcn_9 = 16'b1011001001011101;
    Lcn_10 = 16'b1110000110100010;
    Lcn_11 = 16'b0000011001000111;
    Lcn_12 = 16'b1100111011110011;
    Lcn_13 = 16'b0000101011100010;
    Lcn_14 = 16'b0101100111011001;
    Lcn_15 = 16'b0010000001001110;
    Lcn_16 = 16'b1001110010010110;
    Lcn_17 = 16'b0011001000101110;
    Lcn_18 = 16'b1011001110111011;
    Lcn_19 = 16'b0001011111100100;
    Lcn_20 = 16'b1101010101010010;
    Lcn_21 = 16'b0000110010001110;
    Lcn_22 = 16'b0100001000100101;
    Lcn_23 = 16'b1010001000000001;
    Lcn_24 = 16'b1110000001001000;
    Lcn_25 = 16'b0011100111010110;
    Lcn_26 = 16'b1101001000101011;
    Lcn_27 = 16'b1001011011101110;
    Lcn_28 = 16'b1100000010101010;
    Lcn_29 = 16'b0111011010011001;
    Lcn_30 = 16'b1110101110011001;
    Lcn_31 = 16'b0011000101000111;
    
    #20;
    Lcn_0 = 16'b0111011001110110;
    Lcn_1 = 16'b0001100111011100;
    Lcn_2 = 16'b1101000100110110;
    Lcn_3 = 16'b0010110111110110;
    Lcn_4 = 16'b0110101011110001;
    Lcn_5 = 16'b1001000000000000;
    Lcn_6 = 16'b0110110010010010;
    Lcn_7 = 16'b1100110101101010;
    Lcn_8 = 16'b1001011111101100;
    Lcn_9 = 16'b0011111001011011;
    Lcn_10 = 16'b0100011001101101;
    Lcn_11 = 16'b1011110111110000;
    Lcn_12 = 16'b0100001010011100;
    Lcn_13 = 16'b1000011101100001;
    Lcn_14 = 16'b1111110110001010;
    Lcn_15 = 16'b0011111111010110;
    Lcn_16 = 16'b1010101011100001;
    Lcn_17 = 16'b1100001101011111;
    Lcn_18 = 16'b0010011010111010;
    Lcn_19 = 16'b1000011101101000;
    Lcn_20 = 16'b1010100101101101;
    Lcn_21 = 16'b1010110010101001;
    Lcn_22 = 16'b0101101101010100;
    Lcn_23 = 16'b1111001000101100;
    Lcn_24 = 16'b1110100111010000;
    Lcn_25 = 16'b1100100110000110;
    Lcn_26 = 16'b1010110111010000;
    Lcn_27 = 16'b1101110101101001;
    Lcn_28 = 16'b1101101111101000;
    Lcn_29 = 16'b0100011010001111;
    Lcn_30 = 16'b0011011100110000;
    Lcn_31 = 16'b0010010110111100;
    
    #20;
    Lcn_0 = 16'b0010001101101000;
    Lcn_1 = 16'b1000111010110110;
    Lcn_2 = 16'b0101110101111111;
    Lcn_3 = 16'b0100010010111101;
    Lcn_4 = 16'b0111001111101010;
    Lcn_5 = 16'b1110111001111001;
    Lcn_6 = 16'b0010100001010111;
    Lcn_7 = 16'b0100100110010100;
    Lcn_8 = 16'b0000010110011101;
    Lcn_9 = 16'b1001001000110011;
    Lcn_10 = 16'b0010001011111100;
    Lcn_11 = 16'b1000000101100111;
    Lcn_12 = 16'b1000010110010110;
    Lcn_13 = 16'b0101011011000101;
    Lcn_14 = 16'b0010111111111101;
    Lcn_15 = 16'b1111111111001010;
    Lcn_16 = 16'b0100001001011110;
    Lcn_17 = 16'b0001000110011000;
    Lcn_18 = 16'b0110001011000000;
    Lcn_19 = 16'b0111011111001001;
    Lcn_20 = 16'b0001101000010001;
    Lcn_21 = 16'b1001010111011111;
    Lcn_22 = 16'b0111011010100001;
    Lcn_23 = 16'b0011000011111100;
    Lcn_24 = 16'b0010100000010000;
    Lcn_25 = 16'b1011000001011011;
    Lcn_26 = 16'b1100011001011111;
    Lcn_27 = 16'b0110100001111101;
    Lcn_28 = 16'b1110001110010100;
    Lcn_29 = 16'b0000000001000010;
    Lcn_30 = 16'b1011101010010100;
    Lcn_31 = 16'b1011101100010110;
    
    #20;
    Lcn_0 = 16'b0110101111000111;
    Lcn_1 = 16'b1101001000010100;
    Lcn_2 = 16'b0000110011110010;
    Lcn_3 = 16'b0000000010101100;
    Lcn_4 = 16'b0001001010010101;
    Lcn_5 = 16'b1011101110110011;
    Lcn_6 = 16'b1011011101000001;
    Lcn_7 = 16'b0111000100110011;
    Lcn_8 = 16'b0101110000110101;
    Lcn_9 = 16'b1010011111001101;
    Lcn_10 = 16'b0101110110001001;
    Lcn_11 = 16'b0100101001100100;
    Lcn_12 = 16'b1110101010000100;
    Lcn_13 = 16'b1111010000101011;
    Lcn_14 = 16'b1110100101000101;
    Lcn_15 = 16'b1100100100011010;
    Lcn_16 = 16'b0111011011010111;
    Lcn_17 = 16'b1100011100001010;
    Lcn_18 = 16'b1011001000100110;
    Lcn_19 = 16'b1001010010110111;
    Lcn_20 = 16'b1001101000010110;
    Lcn_21 = 16'b0011100001100100;
    Lcn_22 = 16'b1010010011111010;
    Lcn_23 = 16'b0110110001011010;
    Lcn_24 = 16'b0010010001011000;
    Lcn_25 = 16'b0000111001100110;
    Lcn_26 = 16'b0011111110001011;
    Lcn_27 = 16'b0001110001011111;
    Lcn_28 = 16'b0110001001110011;
    Lcn_29 = 16'b0011001100100000;
    Lcn_30 = 16'b1110111111101101;
    Lcn_31 = 16'b1011000001101111;
    
    #20;
    Lcn_0 = 16'b0010110100100110;
    Lcn_1 = 16'b0000010111111101;
    Lcn_2 = 16'b1101010111000000;
    Lcn_3 = 16'b0101100100100010;
    Lcn_4 = 16'b1110100001101001;
    Lcn_5 = 16'b0010000000100011;
    Lcn_6 = 16'b1000011011101010;
    Lcn_7 = 16'b0000000001010010;
    Lcn_8 = 16'b0101101110011100;
    Lcn_9 = 16'b1100111101001101;
    Lcn_10 = 16'b0010000101011000;
    Lcn_11 = 16'b1011101111111000;
    Lcn_12 = 16'b0111110000110001;
    Lcn_13 = 16'b0111111000110000;
    Lcn_14 = 16'b0100101101101000;
    Lcn_15 = 16'b1100110111001010;
    Lcn_16 = 16'b1101011111101110;
    Lcn_17 = 16'b1111011011010100;
    Lcn_18 = 16'b0010011101010110;
    Lcn_19 = 16'b1011100001100101;
    Lcn_20 = 16'b1001101100110111;
    Lcn_21 = 16'b0001101111001111;
    Lcn_22 = 16'b0100011100001011;
    Lcn_23 = 16'b1011011000100010;
    Lcn_24 = 16'b0001000010110100;
    Lcn_25 = 16'b1101001101010100;
    Lcn_26 = 16'b1010000000100011;
    Lcn_27 = 16'b0010110011011011;
    Lcn_28 = 16'b1100100110001100;
    Lcn_29 = 16'b1011000010000011;
    Lcn_30 = 16'b1001000010011010;
    Lcn_31 = 16'b1111100111011100;
    
    #20;
    Lcn_0 = 16'b1000110101110100;
    Lcn_1 = 16'b0010100001011101;
    Lcn_2 = 16'b1111100111100001;
    Lcn_3 = 16'b0101111101100100;
    Lcn_4 = 16'b1011111011000001;
    Lcn_5 = 16'b0000011101010000;
    Lcn_6 = 16'b1001111000101010;
    Lcn_7 = 16'b1101000110011010;
    Lcn_8 = 16'b1100011000000110;
    Lcn_9 = 16'b0101011110001001;
    Lcn_10 = 16'b0111100011011011;
    Lcn_11 = 16'b0100001011011001;
    Lcn_12 = 16'b0001100110100010;
    Lcn_13 = 16'b1000100010010101;
    Lcn_14 = 16'b0011110011011101;
    Lcn_15 = 16'b0001110111111101;
    Lcn_16 = 16'b1111100100001010;
    Lcn_17 = 16'b0000001000000100;
    Lcn_18 = 16'b0110110011101001;
    Lcn_19 = 16'b1010011110110001;
    Lcn_20 = 16'b0010000100000011;
    Lcn_21 = 16'b1111101101010011;
    Lcn_22 = 16'b1101111001000100;
    Lcn_23 = 16'b0000011000101010;
    Lcn_24 = 16'b1111110011000010;
    Lcn_25 = 16'b1101100001110000;
    Lcn_26 = 16'b0011100000111110;
    Lcn_27 = 16'b0110111101101100;
    Lcn_28 = 16'b0110101000000111;
    Lcn_29 = 16'b1001111010101011;
    Lcn_30 = 16'b0010110000100011;
    Lcn_31 = 16'b0001110000011000;
    
    #20;
    Lcn_0 = 16'b0011101000001001;
    Lcn_1 = 16'b0010101011110011;
    Lcn_2 = 16'b1111101111000011;
    Lcn_3 = 16'b1111011101101000;
    Lcn_4 = 16'b1001111010110100;
    Lcn_5 = 16'b0000011101100100;
    Lcn_6 = 16'b1110110101101100;
    Lcn_7 = 16'b0001100100000010;
    Lcn_8 = 16'b0010100111001101;
    Lcn_9 = 16'b1010110111110000;
    Lcn_10 = 16'b1111100101100011;
    Lcn_11 = 16'b0101100111110100;
    Lcn_12 = 16'b1111000010110110;
    Lcn_13 = 16'b1101110111010111;
    Lcn_14 = 16'b1010000100010111;
    Lcn_15 = 16'b0100100110011011;
    Lcn_16 = 16'b0110011111000010;
    Lcn_17 = 16'b0101100011111100;
    Lcn_18 = 16'b1101110011100001;
    Lcn_19 = 16'b0010101011000010;
    Lcn_20 = 16'b0011010111100101;
    Lcn_21 = 16'b0100100110101001;
    Lcn_22 = 16'b1111010001110111;
    Lcn_23 = 16'b1101110000111101;
    Lcn_24 = 16'b1111010010111011;
    Lcn_25 = 16'b0101110010101111;
    Lcn_26 = 16'b1110100110000110;
    Lcn_27 = 16'b1001001001001001;
    Lcn_28 = 16'b1110100100110100;
    Lcn_29 = 16'b1010000110000110;
    Lcn_30 = 16'b0001001110110110;
    Lcn_31 = 16'b0100111100011010;
    
    #20;
    Lcn_0 = 16'b0011011100011000;
    Lcn_1 = 16'b1110100010010100;
    Lcn_2 = 16'b0100110101010100;
    Lcn_3 = 16'b1111100100101010;
    Lcn_4 = 16'b1110100000100110;
    Lcn_5 = 16'b1011010100000001;
    Lcn_6 = 16'b0110100010001001;
    Lcn_7 = 16'b1101000000010111;
    Lcn_8 = 16'b0011110111000000;
    Lcn_9 = 16'b1010101111101100;
    Lcn_10 = 16'b1100000001110000;
    Lcn_11 = 16'b0111000110011101;
    Lcn_12 = 16'b1000110110111011;
    Lcn_13 = 16'b1001011010000100;
    Lcn_14 = 16'b1000010011111000;
    Lcn_15 = 16'b0011101001000010;
    Lcn_16 = 16'b0101011010101110;
    Lcn_17 = 16'b1000001110100011;
    Lcn_18 = 16'b1110001110101101;
    Lcn_19 = 16'b0101100101000001;
    Lcn_20 = 16'b0110101010011100;
    Lcn_21 = 16'b1001011101101101;
    Lcn_22 = 16'b0011110001110010;
    Lcn_23 = 16'b1011000010111000;
    Lcn_24 = 16'b1000100011010010;
    Lcn_25 = 16'b1101000011000011;
    Lcn_26 = 16'b1011010100111110;
    Lcn_27 = 16'b1101110110100011;
    Lcn_28 = 16'b1111100001100000;
    Lcn_29 = 16'b0001110010110100;
    Lcn_30 = 16'b1011011100001110;
    Lcn_31 = 16'b1110100011011000;
    
    #20;
    Lcn_0 = 16'b1001011101101000;
    Lcn_1 = 16'b0110000111111000;
    Lcn_2 = 16'b0011101001100011;
    Lcn_3 = 16'b0001000111000100;
    Lcn_4 = 16'b0001011110011101;
    Lcn_5 = 16'b1110010111100011;
    Lcn_6 = 16'b1001011010010001;
    Lcn_7 = 16'b0101010100101101;
    Lcn_8 = 16'b1111101010110011;
    Lcn_9 = 16'b0010011100010111;
    Lcn_10 = 16'b1100011001010100;
    Lcn_11 = 16'b1010101001100100;
    Lcn_12 = 16'b1010101011101000;
    Lcn_13 = 16'b1111001110100010;
    Lcn_14 = 16'b1100110010100000;
    Lcn_15 = 16'b0110001000011111;
    Lcn_16 = 16'b0011100010110000;
    Lcn_17 = 16'b0100110000100010;
    Lcn_18 = 16'b1110010101010000;
    Lcn_19 = 16'b1011001111101011;
    Lcn_20 = 16'b1110010011101110;
    Lcn_21 = 16'b0110101110101010;
    Lcn_22 = 16'b1111111100111001;
    Lcn_23 = 16'b0111000100110011;
    Lcn_24 = 16'b1111001000101111;
    Lcn_25 = 16'b1000000011000000;
    Lcn_26 = 16'b0101111000011100;
    Lcn_27 = 16'b1000111011000101;
    Lcn_28 = 16'b0111010111010111;
    Lcn_29 = 16'b0000100010011100;
    Lcn_30 = 16'b0010111010111001;
    Lcn_31 = 16'b1001011110111010;
    
    #20;
    Lcn_0 = 16'b0101011010101110;
    Lcn_1 = 16'b0110011110000101;
    Lcn_2 = 16'b0101010101101100;
    Lcn_3 = 16'b1001100011101011;
    Lcn_4 = 16'b0101100011111010;
    Lcn_5 = 16'b1001001000101100;
    Lcn_6 = 16'b0000010110001001;
    Lcn_7 = 16'b1101100101010101;
    Lcn_8 = 16'b0001110010010110;
    Lcn_9 = 16'b1000110001110111;
    Lcn_10 = 16'b1011010010010001;
    Lcn_11 = 16'b1000011111100000;
    Lcn_12 = 16'b1100011000100010;
    Lcn_13 = 16'b0101110010110000;
    Lcn_14 = 16'b0111000110010000;
    Lcn_15 = 16'b1111010110110010;
    Lcn_16 = 16'b1111001010011101;
    Lcn_17 = 16'b0100000110101111;
    Lcn_18 = 16'b0110000110111011;
    Lcn_19 = 16'b1000100011000011;
    Lcn_20 = 16'b0110010010000000;
    Lcn_21 = 16'b0010101010001111;
    Lcn_22 = 16'b0010010000110011;
    Lcn_23 = 16'b0111110110110111;
    Lcn_24 = 16'b0101001001011010;
    Lcn_25 = 16'b0101000100011001;
    Lcn_26 = 16'b0110100011110101;
    Lcn_27 = 16'b1111010011000100;
    Lcn_28 = 16'b0111101010000110;
    Lcn_29 = 16'b0101001111110110;
    Lcn_30 = 16'b1010110101001100;
    Lcn_31 = 16'b1010111000000011;
    
    #20;
    Lcn_0 = 16'b0011111100100010;
    Lcn_1 = 16'b0111111101110100;
    Lcn_2 = 16'b1111110101011000;
    Lcn_3 = 16'b0101001010111111;
    Lcn_4 = 16'b1101100111000101;
    Lcn_5 = 16'b1111000110100011;
    Lcn_6 = 16'b0001101011000010;
    Lcn_7 = 16'b0001000110010001;
    Lcn_8 = 16'b0101110001010111;
    Lcn_9 = 16'b1010100111111011;
    Lcn_10 = 16'b1000111001101010;
    Lcn_11 = 16'b1000100100110101;
    Lcn_12 = 16'b0101111111100100;
    Lcn_13 = 16'b1110111001000000;
    Lcn_14 = 16'b1100000010000100;
    Lcn_15 = 16'b0101111000000011;
    Lcn_16 = 16'b1100011111111001;
    Lcn_17 = 16'b0010101111001011;
    Lcn_18 = 16'b0011111011010010;
    Lcn_19 = 16'b0001000000101001;
    Lcn_20 = 16'b0110011010000100;
    Lcn_21 = 16'b0110111000100010;
    Lcn_22 = 16'b0010100011001111;
    Lcn_23 = 16'b1101000100111000;
    Lcn_24 = 16'b0001010000101110;
    Lcn_25 = 16'b0101111000011011;
    Lcn_26 = 16'b1100101101011001;
    Lcn_27 = 16'b0010111011010111;
    Lcn_28 = 16'b0111011000110000;
    Lcn_29 = 16'b0100011100011000;
    Lcn_30 = 16'b0001100100101011;
    Lcn_31 = 16'b1110110010001100;
    
    #20;
    Lcn_0 = 16'b0011111110101110;
    Lcn_1 = 16'b0011101101011000;
    Lcn_2 = 16'b1011101110001101;
    Lcn_3 = 16'b0000011110101001;
    Lcn_4 = 16'b1011101100001110;
    Lcn_5 = 16'b1011111111110100;
    Lcn_6 = 16'b1001100000010001;
    Lcn_7 = 16'b0110101100001000;
    Lcn_8 = 16'b1010100111111101;
    Lcn_9 = 16'b0111000100101100;
    Lcn_10 = 16'b0010101011010010;
    Lcn_11 = 16'b0011011101110010;
    Lcn_12 = 16'b0000101111100001;
    Lcn_13 = 16'b1011001100000001;
    Lcn_14 = 16'b1100010001101010;
    Lcn_15 = 16'b0101100100000101;
    Lcn_16 = 16'b0000011010111101;
    Lcn_17 = 16'b0011101001110101;
    Lcn_18 = 16'b0011110010100100;
    Lcn_19 = 16'b1010011110110001;
    Lcn_20 = 16'b0101111100000000;
    Lcn_21 = 16'b0010100011001111;
    Lcn_22 = 16'b0001010111101001;
    Lcn_23 = 16'b1000010011000101;
    Lcn_24 = 16'b0111111110001110;
    Lcn_25 = 16'b0011100011100100;
    Lcn_26 = 16'b0101010010000000;
    Lcn_27 = 16'b1011001011100110;
    Lcn_28 = 16'b1101010101010011;
    Lcn_29 = 16'b1000110100111111;
    Lcn_30 = 16'b0101010001001101;
    Lcn_31 = 16'b0010110101000110;
    
    #20;
    Lcn_0 = 16'b0110010011001011;
    Lcn_1 = 16'b1010101011011011;
    Lcn_2 = 16'b1100001001101001;
    Lcn_3 = 16'b0101101110010011;
    Lcn_4 = 16'b0000001101100111;
    Lcn_5 = 16'b0011101010010110;
    Lcn_6 = 16'b0111011010101010;
    Lcn_7 = 16'b0011000000111011;
    Lcn_8 = 16'b1100011001111101;
    Lcn_9 = 16'b0000100101011011;
    Lcn_10 = 16'b0100110110000101;
    Lcn_11 = 16'b0010010000001010;
    Lcn_12 = 16'b0110111001111000;
    Lcn_13 = 16'b1100100010111000;
    Lcn_14 = 16'b1111111001011011;
    Lcn_15 = 16'b1001111011010110;
    Lcn_16 = 16'b0011100000000010;
    Lcn_17 = 16'b1000101011111011;
    Lcn_18 = 16'b1101000111000001;
    Lcn_19 = 16'b0110000110001101;
    Lcn_20 = 16'b0011100010001010;
    Lcn_21 = 16'b1011110101011000;
    Lcn_22 = 16'b0001100010101110;
    Lcn_23 = 16'b1001010001001001;
    Lcn_24 = 16'b1000110101111000;
    Lcn_25 = 16'b0110001001000011;
    Lcn_26 = 16'b0110101001000100;
    Lcn_27 = 16'b1110100110110011;
    Lcn_28 = 16'b0101101101111111;
    Lcn_29 = 16'b1010100000001101;
    Lcn_30 = 16'b1101110000001100;
    Lcn_31 = 16'b1101101000000011;
    
    #20;
    Lcn_0 = 16'b0000001101001111;
    Lcn_1 = 16'b1000100110010101;
    Lcn_2 = 16'b1101001001100000;
    Lcn_3 = 16'b1100111100000110;
    Lcn_4 = 16'b0100000110100100;
    Lcn_5 = 16'b1011010000011011;
    Lcn_6 = 16'b1100000111101000;
    Lcn_7 = 16'b0000000111001111;
    Lcn_8 = 16'b0000100111111010;
    Lcn_9 = 16'b0011101100011111;
    Lcn_10 = 16'b1010111100011001;
    Lcn_11 = 16'b1111001010110110;
    Lcn_12 = 16'b0000100100001101;
    Lcn_13 = 16'b1011111010010111;
    Lcn_14 = 16'b1111111111100011;
    Lcn_15 = 16'b0100111001011000;
    Lcn_16 = 16'b0100100010101111;
    Lcn_17 = 16'b1011100100001011;
    Lcn_18 = 16'b1100011101111011;
    Lcn_19 = 16'b0101101000100110;
    Lcn_20 = 16'b0011110111000001;
    Lcn_21 = 16'b1010111110001001;
    Lcn_22 = 16'b1101001100001101;
    Lcn_23 = 16'b0000110110100001;
    Lcn_24 = 16'b0000111110001111;
    Lcn_25 = 16'b1001100100011011;
    Lcn_26 = 16'b1010111110111011;
    Lcn_27 = 16'b0010100001110011;
    Lcn_28 = 16'b1111111000110011;
    Lcn_29 = 16'b0111010111111000;
    Lcn_30 = 16'b0011100110010100;
    Lcn_31 = 16'b1110000101100000;
    
    #20;
    Lcn_0 = 16'b0101011011011100;
    Lcn_1 = 16'b1011101100111001;
    Lcn_2 = 16'b1110101011101011;
    Lcn_3 = 16'b0010001111100100;
    Lcn_4 = 16'b1011001110101100;
    Lcn_5 = 16'b1011011101011111;
    Lcn_6 = 16'b0111111011001010;
    Lcn_7 = 16'b0100111010110010;
    Lcn_8 = 16'b0000011110110100;
    Lcn_9 = 16'b0011110000011100;
    Lcn_10 = 16'b1000100100101101;
    Lcn_11 = 16'b0011110111011000;
    Lcn_12 = 16'b1010000110010101;
    Lcn_13 = 16'b1010010100100101;
    Lcn_14 = 16'b0010001001010101;
    Lcn_15 = 16'b1111110101101000;
    Lcn_16 = 16'b1110011100010011;
    Lcn_17 = 16'b0010101111111010;
    Lcn_18 = 16'b0101110101000011;
    Lcn_19 = 16'b1101101001001000;
    Lcn_20 = 16'b0010111101011010;
    Lcn_21 = 16'b1101111010110000;
    Lcn_22 = 16'b1010001001000011;
    Lcn_23 = 16'b1001100010101011;
    Lcn_24 = 16'b1000100110001010;
    Lcn_25 = 16'b1111100001100110;
    Lcn_26 = 16'b0111101101100011;
    Lcn_27 = 16'b0011011000101110;
    Lcn_28 = 16'b1100001111001100;
    Lcn_29 = 16'b0100011001000101;
    Lcn_30 = 16'b0001001101110010;
    Lcn_31 = 16'b1101001101111100;
    
    #20;
    Lcn_0 = 16'b0101010100100110;
    Lcn_1 = 16'b0111011111111100;
    Lcn_2 = 16'b1100000101110010;
    Lcn_3 = 16'b0011001010011110;
    Lcn_4 = 16'b0110101100101100;
    Lcn_5 = 16'b0111000001010110;
    Lcn_6 = 16'b0100010100010010;
    Lcn_7 = 16'b0101001100010111;
    Lcn_8 = 16'b1111100100111010;
    Lcn_9 = 16'b0100111100011010;
    Lcn_10 = 16'b1111101000111101;
    Lcn_11 = 16'b0000000110011010;
    Lcn_12 = 16'b1111100010010011;
    Lcn_13 = 16'b0111010100000011;
    Lcn_14 = 16'b1011110101010010;
    Lcn_15 = 16'b0001111101010110;
    Lcn_16 = 16'b0011011110101011;
    Lcn_17 = 16'b1100011000011010;
    Lcn_18 = 16'b0000011011001000;
    Lcn_19 = 16'b0110001011110011;
    Lcn_20 = 16'b0110010010010101;
    Lcn_21 = 16'b1010100101100000;
    Lcn_22 = 16'b0100110111100000;
    Lcn_23 = 16'b1000111100011011;
    Lcn_24 = 16'b0111100001000000;
    Lcn_25 = 16'b0011011000010100;
    Lcn_26 = 16'b0011111001111011;
    Lcn_27 = 16'b1100111010100110;
    Lcn_28 = 16'b1110100101000000;
    Lcn_29 = 16'b1010000011110001;
    Lcn_30 = 16'b1011101101100100;
    Lcn_31 = 16'b1001110110100001;
    
    #20;
    Lcn_0 = 16'b0101000000110100;
    Lcn_1 = 16'b0011011101010100;
    Lcn_2 = 16'b1110011100101100;
    Lcn_3 = 16'b0101011110110010;
    Lcn_4 = 16'b1000000111110111;
    Lcn_5 = 16'b0011011101111001;
    Lcn_6 = 16'b1111110100011010;
    Lcn_7 = 16'b0100110000010100;
    Lcn_8 = 16'b1010011011000011;
    Lcn_9 = 16'b0111000001101101;
    Lcn_10 = 16'b1000111101110000;
    Lcn_11 = 16'b0000110011000101;
    Lcn_12 = 16'b1100011010111000;
    Lcn_13 = 16'b1010001011111100;
    Lcn_14 = 16'b1000100101101111;
    Lcn_15 = 16'b1111100000110100;
    Lcn_16 = 16'b1000100100010100;
    Lcn_17 = 16'b0100100111100001;
    Lcn_18 = 16'b1110111010010001;
    Lcn_19 = 16'b1101011100000110;
    Lcn_20 = 16'b0111001110100010;
    Lcn_21 = 16'b1011001001001111;
    Lcn_22 = 16'b0000001100000101;
    Lcn_23 = 16'b0111100110000010;
    Lcn_24 = 16'b1100011011001000;
    Lcn_25 = 16'b0111100111000000;
    Lcn_26 = 16'b1011001010101010;
    Lcn_27 = 16'b1110100011100011;
    Lcn_28 = 16'b0110111100111000;
    Lcn_29 = 16'b0110011110001000;
    Lcn_30 = 16'b0011010000100100;
    Lcn_31 = 16'b1111011100001000;
    
    #20;
    Lcn_0 = 16'b0110100110100100;
    Lcn_1 = 16'b1110110000000000;
    Lcn_2 = 16'b0111111001000111;
    Lcn_3 = 16'b0011011010010101;
    Lcn_4 = 16'b0010010010111111;
    Lcn_5 = 16'b0010011010001110;
    Lcn_6 = 16'b0100000010010001;
    Lcn_7 = 16'b0111001101011111;
    Lcn_8 = 16'b1110010101111101;
    Lcn_9 = 16'b1011011110010111;
    Lcn_10 = 16'b1101111011011010;
    Lcn_11 = 16'b0111001101000101;
    Lcn_12 = 16'b1101010001011111;
    Lcn_13 = 16'b0010011111101101;
    Lcn_14 = 16'b0001101110101111;
    Lcn_15 = 16'b0110010001000111;
    Lcn_16 = 16'b1101111110011111;
    Lcn_17 = 16'b1010011011011111;
    Lcn_18 = 16'b0100000111101100;
    Lcn_19 = 16'b0101010010111110;
    Lcn_20 = 16'b0100011010011101;
    Lcn_21 = 16'b0011110001101000;
    Lcn_22 = 16'b1011111111110100;
    Lcn_23 = 16'b1111110110011010;
    Lcn_24 = 16'b0111100011111010;
    Lcn_25 = 16'b0110110110001010;
    Lcn_26 = 16'b1011010101110101;
    Lcn_27 = 16'b0110010010111110;
    Lcn_28 = 16'b0011001101010010;
    Lcn_29 = 16'b1110011110000010;
    Lcn_30 = 16'b0000101010010011;
    Lcn_31 = 16'b0100001101101000;
    
    #20;
    Lcn_0 = 16'b1010010110010011;
    Lcn_1 = 16'b1111101111100011;
    Lcn_2 = 16'b0100000001011001;
    Lcn_3 = 16'b1111110010110011;
    Lcn_4 = 16'b0100000000000010;
    Lcn_5 = 16'b1100110111101010;
    Lcn_6 = 16'b0111001010001100;
    Lcn_7 = 16'b1001111110100110;
    Lcn_8 = 16'b0011001011101011;
    Lcn_9 = 16'b0111000001011001;
    Lcn_10 = 16'b0110010101000000;
    Lcn_11 = 16'b1100001110101110;
    Lcn_12 = 16'b1100101011001111;
    Lcn_13 = 16'b1110101110100111;
    Lcn_14 = 16'b0101101010011010;
    Lcn_15 = 16'b0010100000101010;
    Lcn_16 = 16'b1100011001100110;
    Lcn_17 = 16'b0000000010001000;
    Lcn_18 = 16'b1100101111111100;
    Lcn_19 = 16'b0010010111110000;
    Lcn_20 = 16'b1111000010000110;
    Lcn_21 = 16'b1001010010111101;
    Lcn_22 = 16'b1101011001001011;
    Lcn_23 = 16'b1000111000111001;
    Lcn_24 = 16'b0001110110011010;
    Lcn_25 = 16'b0000001110010001;
    Lcn_26 = 16'b1111010110100000;
    Lcn_27 = 16'b1101000001010110;
    Lcn_28 = 16'b0000001111110000;
    Lcn_29 = 16'b1000111001011111;
    Lcn_30 = 16'b1101111101001000;
    Lcn_31 = 16'b1111101011101000;
    #90;

    $stop;
end



endmodule

